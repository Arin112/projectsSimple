﻿module vReg16
/*
далее представлен 16-ти разрядный регистр
когда бит load равен единице происходит параллельная загрузка из data
когда бит load равен нулю происходит последовательная загрузка из бита b
*/
(
	input [15:0] data,
	input b,
	input load, clk,
	output reg [15:0] q // ключевое слово reg показывает, что под q будет выделено место
); // reg переменные можно менять по возникновению событий

	always @ (posedge clk) // дословно - вызывать последующий блок begin ... end всегда, когда сигнал clk менят значение с нуля на единицу
	// posedge - positive edge - положительный фронт
	// аналогично существует событие negedge
	// также события можно назначать на изменение любого из входных сигналов при помощи always @*
	// на изменение нескольких сигналов always @(a or b or c)
	begin
		if (load)
			q <= data; // <= - неблокирующее присваивание - каждая строчка с <= будет выполнена параллельно
		else begin
			q = q >> 1; // сдвиг регистра
			// тут присваивание блокирующее - строки будут выполнены 'последовательно'
			// в кавычках так как в действительности всё произойдёт за 1 такт
			q[15] = b;
		end
	end

endmodule
