﻿module sum4
(
input [3:0] a, // четырёхбитное число
input [3:0] b, // или же массив из четырех бит, что то же самое
input cin,
output [3:0] c, // ответ
output cout
);
wire [3:0] couts; // wire это 'тип данных' означающий,
// что внутри схемы не будует создаваться отдельных регистров или ячеек для хранения,
// а все использования таких переменных будут заменены на их значения
// в wire возможно использовать только непрерывное присваивание
// все входные input сигналы - wire
vSum inst0(.a(a[0]), .b(b[0]), .cin(cin), .c(c[0]), .cout(couts[0]));
// так в verilog используются модули - в данном случа ранее написанный vSum
// имя_модуля имя_экземпляра(.имя_входного_сигнала(имя), .имя_выходного_сигнала(имя));
// при создании inst0 была создана непрерывная цепочка соединяющая a[0], b[0], cin и c[0], couts[0]
genvar x; // специальная переменная, которую можно использовать для итерации внутри генератора
generate // специальный блок, внутри которого можно создавать множество экземпляров модуля
	for(x = 1; x < 4; x = x + 1)begin : _gen1
		// практически обычный цикл в стиле Си, разве что поле begin стоит двоеточие,
		// а после него название цикла(любое, тут все циклы именные)
		vSum insts(.a(a[x]), .b(b[x]), .c(c[x]), .cin(couts[x-1]), .cout(couts[x]));
	end
endgenerate
assign cout = couts[3]; // бит переноса последней суммы это бит переноса этого модуля

endmodule
