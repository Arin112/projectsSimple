module ALU
(
	input [7:0] a,b,  	// два восьмибитных входа                 
	input [3:0] op,		// индекс операции
	output reg [7:0] res, 	// результат операции
	// ключевое слово reg означает, что под переменную будет выделена память в блоке
	// по умолчанию тип wire
	output cout 		// флаг переполнения
);

	wire [8:0] tmp;
	// wire - тип данных, означающий, что переменная не будет существовать как ячейка памяти в блоке
	// дословно - провод, что очень точно отражает суть происходящего
	// провода как бы висят в воздухе - не занимают места, только логические вентили

	assign cout = tmp[8];
	// так провода соединяют - теперь cout имеет точно такое же значени что и восьмой бит tmp

	assign tmp = {1'b0,a} + {1'b0,b};
	// фигурные скобки объединяют перечисленные в них переменные
	// в первом случае нулевой бит и wire переменную a
	// во втором то же самое с b
	// операция + это обычное сложение
	// вся замысловатая конструкция выше нужна для того чтобы присвоить в cout бит,
	// который всегда будет означать будет ли переполнение при сложении заданных чисел a и b
	
	always @(*) begin
	// конструкция always @(*) дословно говорит "исполнять последующий блок begin ... end
	// каждый раз, когда какой либо входной сигнал изменит значение"
	
	// case в этом языке похож на switch из других языков, с тем отличием, что одной метке
	// сопоставляется только последующий блок, который либо представляет собой begin ... end
	// либо выражение, заканчивающиеся точкой с запятой
		case(op)
			4'h0: // сложение
				res = a + b ; 
			4'h1: // вычитание
				res = a - b ;
			4'h2: // умножение
				res = a * b;
			4'h3: // деление
				res = a/b;
			4'h4: // побитовый сдвиг влево на 1 бит
				res = a<<1;
			4'h5: // побитовый сдвиг вправо на 1 бит
				res = a>>1;
			4'h6: // циклический сдвиг влево
				res = {a[6:0],a[7]};
			4'h7: // циклический сдвиг вправо
				res = {a[0],a[7:1]};
			4'h8: //  побитовое и
				res = a & b;
			4'h9: //  побитовое или
				res = a | b;
			4'hA: //  побитовое исключающее или 
				res = a ^ b;
			4'hB: //  побитовое отрицание побитового исключающего или
				res = ~(a | b);
			4'hC: // побитовое отрицание побитового и
				res = ~(a & b);
			4'hD: // побитовое отрцание побитового исключающего и
				res = ~(a ^ b);
			4'hE: // сравнение больше чем
				res = (a>b)?8'd1:8'd0 ;
			4'hF: // сравнение меньше чем
				res = (a==b)?8'd1:8'd0 ;
			default: res = a + b ; // не должно быть выполнено никогда, кроме отладочных высокоимпедентных состояний
			// высокоимпедентное состояние - третье состояние в котором может находиться бит
			// возможно только в симуляции для отладки, не может быть синтезировано в микросхеме
		endcase
	end

endmodule
