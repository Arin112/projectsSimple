﻿module vSum // модуль складывает два бита с использованием битов переноса
// вообще говоря, в verilog сложение шеснадцатибитных чисел можно написать как a + b
// но написание сумматора это хорошая возможность продемонстрировать основы языка
(
input a, // первое слагаемое
input b, // второе слагаемое
input cin, // бит переноса с предыдущего слагаемого
output c, // сумма
output cout // бит переноса на следующее слагаемое
);
// здесь возможно только непрерывное присваивание (в глобальной области)
// в действительности это не приваивание в привычном смысле
assign c = a ^ b ^ cin; // нахождение суммы
// неверное прочтение записи выше - 'положить в ячейку c значение выражения a^b^cin над переменными a, b и cin'
// правильное прочтение - 'сконфигурировать логические вентили таким образом, что выходной сигнал c будет равен выражению a^b^cin над входными сигналами a, b и cin'
// таким образом становится понятно, что в данном случае выстраивается непрерывная цепочка из логических вентелей соединяющая входные и выходные сигналы
assign cout = (a & b) || (a & cin) || (b & cin); // бит переноса
// результат непрерывного присваивания меняется как только меняются входные сигналы
endmodule
